module flags();

endmodule